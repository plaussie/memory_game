`ifndef _game_params
`define _game_params

//Colors
`define BACKGROUND_TXT_COLOR 12'hf_8_b
`define BACKGROUND_COLOR 12'h8_8_f
`define BUTTON_TXT_COLOR 12'h8_8_f
`define BUTTON_COLOR 12'hf_8_b

//Start Button Params
`define START_BUTTON_X_POS 412
`define START_BUTTON_Y_POS 328
`define START_BUTTON_WIDTH 200
`define START_BUTTON_HEIGHT 112
`define START_BUTTON_ROM_WIDTH_SIZE 8
`define START_BUTTON_ROM_HEIGHT_SIZE 8
`define START_BUTTON_ROM_PATH "start_button.data"

//Options Button Params
`define OPTIONS_BUTTON_X_POS 106
`define OPTIONS_BUTTON_Y_POS 328
`define OPTIONS_BUTTON_WIDTH 200
`define OPTIONS_BUTTON_HEIGHT 112
`define OPTIONS_BUTTON_ROM_WIDTH_SIZE 8
`define OPTIONS_BUTTON_ROM_HEIGHT_SIZE 8
`define OPTIONS_BUTTON_ROM_PATH "options_button.data"

//Easy Button Params
`define EASY_BUTTON_X_POS 106
`define EASY_BUTTON_Y_POS 328
`define EASY_BUTTON_WIDTH 200
`define EASY_BUTTON_HEIGHT 112
`define EASY_BUTTON_ROM_WIDTH_SIZE 8
`define EASY_BUTTON_ROM_HEIGHT_SIZE 8
`define EASY_BUTTON_ROM_PATH "easy_button.data"

//Normal Button Params
`define NORMAL_BUTTON_X_POS 412
`define NORMAL_BUTTON_Y_POS 328
`define NORMAL_BUTTON_WIDTH 200
`define NORMAL_BUTTON_HEIGHT 112
`define NORMAL_BUTTON_ROM_WIDTH_SIZE 8
`define NORMAL_BUTTON_ROM_HEIGHT_SIZE 8
`define NORMAL_BUTTON_ROM_PATH "normal_button.data"

//Hard Button Params
`define HARD_BUTTON_X_POS 718
`define HARD_BUTTON_Y_POS 328
`define HARD_BUTTON_WIDTH 200
`define HARD_BUTTON_HEIGHT 112
`define HARD_BUTTON_ROM_WIDTH_SIZE 8
`define HARD_BUTTON_ROM_HEIGHT_SIZE 8
`define HARD_BUTTON_ROM_PATH "hard_button.data"

//Back Button Params
`define BACK_BUTTON_X_POS 724
`define BACK_BUTTON_Y_POS 556
`define BACK_BUTTON_WIDTH 200
`define BACK_BUTTON_HEIGHT 112
`define BACK_BUTTON_ROM_WIDTH_SIZE 8
`define BACK_BUTTON_ROM_HEIGHT_SIZE 8
`define BACK_BUTTON_ROM_PATH "back_button.data"

`endif