`ifndef _cards_macros
`define _cards_macros

//Difficulty Params
`define CARD_MAX_NUM 16
`define CARD_MAX_NUM_SIZE 5

`define CARD_LEVEL_NUM 3
`define CARD_NUM_EASY 8
`define CARD_NUM_NORMAL 12
`define CARD_NUM_HARD 16

//Cards Params
`define CARD_ADDRESS_SIZE 5
`define CARD_COLOR_SIZE 12
`define CARD_STATE_SIZE 2
`define CARD_DATA_SIZE `CARD_COLOR_SIZE+`CARD_STATE_SIZE
`define CARD_YX_POSITION_SIZE 20
`define FIRST_CARD_INDEX 1

`endif