`ifndef _game_params
`define _game_params

//Start Button Params
`define START_BUTTON_X_POS 412
`define START_BUTTON_Y_POS 328
`define START_BUTTON_WIDTH 200
`define START_BUTTON_HEIGHT 112
`define START_BUTTON_ADDRESS_SIZE 16
`define START_BUTTON_ROM_PIXELS_NUM 65536
`define START_BUTTON_ROM_PATH "start_button.data"

//Options Button Params
`define OPTIONS_BUTTON_X_POS 106
`define OPTIONS_BUTTON_Y_POS 328
`define OPTIONS_BUTTON_WIDTH 200
`define OPTIONS_BUTTON_HEIGHT 112
`define OPTIONS_BUTTON_ADDRESS_SIZE 16
`define OPTIONS_BUTTON_ROM_PIXELS_NUM 65536
`define OPTIONS_BUTTON_ROM_PATH "start_button.data"

//Easy Button Params
`define EASY_BUTTON_X_POS 106
`define EASY_BUTTON_Y_POS 328
`define EASY_BUTTON_WIDTH 200
`define EASY_BUTTON_HEIGHT 112
`define EASY_BUTTON_ADDRESS_SIZE 16
`define EASY_BUTTON_ROM_PIXELS_NUM 65536
`define EASY_BUTTON_ROM_PATH "start_button.data"

//Normal Button Params
`define NORMAL_BUTTON_X_POS 412
`define NORMAL_BUTTON_Y_POS 328
`define NORMAL_BUTTON_WIDTH 200
`define NORMAL_BUTTON_HEIGHT 112
`define NORMAL_BUTTON_ADDRESS_SIZE 16
`define NORMAL_BUTTON_ROM_PIXELS_NUM 65536
`define NORMAL_BUTTON_ROM_PATH "start_button.data"

//Hard Button Params
`define HARD_BUTTON_X_POS 718
`define HARD_BUTTON_Y_POS 328
`define HARD_BUTTON_WIDTH 200
`define HARD_BUTTON_HEIGHT 112
`define HARD_BUTTON_ADDRESS_SIZE 16
`define HARD_BUTTON_ROM_PIXELS_NUM 65536
`define HARD_BUTTON_ROM_PATH "start_button.data"

//Back Button Params
`define BACK_BUTTON_X_POS 724
`define BACK_BUTTON_Y_POS 556
`define BACK_BUTTON_WIDTH 200
`define BACK_BUTTON_HEIGHT 112
`define BACK_BUTTON_ADDRESS_SIZE 16
`define BACK_BUTTON_ROM_PIXELS_NUM 65536
`define BACK_BUTTON_ROM_PATH "start_button.data"

`endif